** Profile: "SCHEMATIC1-SR"  [ C:\Users\sarid\OneDrive\Documents\OpAmp\operational amplifier-pspicefiles\schematic1\sr.sim ] 

** Creating circuit file "SR.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../operational amplifier-pspicefiles/operational amplifier.lib" 
* From [PSPICE NETLIST] section of C:\Users\sarid\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
